// set_associative_cache.sv