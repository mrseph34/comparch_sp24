// set_associative_cache_tb.sv
