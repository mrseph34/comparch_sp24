// tb_direct_mapped_cache.sv
