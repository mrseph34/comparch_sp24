// direct_mapped_cache.sv
